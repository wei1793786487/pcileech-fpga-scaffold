//
// PCILeech FPGA.
//
// PCIe BAR PIO controller.
//
// The PCILeech BAR PIO controller allows for easy user-implementation on top
// of the PCILeech AXIS128 PCIe TLP streaming interface.
// The controller consists of a read engine and a write engine and pluggable
// user-implemented PCIe BAR implementations (found at bottom of the file).
//
// Considerations:
// - The core handles 1 DWORD read + 1 DWORD write per CLK max. If a lot of
//   data is written / read from the TLP streaming interface the core may
//   drop packet silently.
// - The core reads 1 DWORD of data (without byte enable) per CLK.
// - The core writes 1 DWORD of data (with byte enable) per CLK.
// - All user-implemented cores must have the same latency in CLKs for the
//   returned read data or else undefined behavior will take place.
// - 32-bit addresses are passed for read/writes. Larger BARs than 4GB are
//   not supported due to addressing constraints. Lower bits (LSBs) are the
//   BAR offset, Higher bits (MSBs) are the 32-bit base address of the BAR.
// - DO NOT edit read/write engines.
// - DO edit pcileech_tlps128_bar_controller (to swap bar implementations).
// - DO edit the bar implementations (at bottom of the file, if neccessary).
//
// Example implementations exists below, swap out any of the example cores
// against a core of your use case, or modify existing cores.
// Following test cores exist (see below in this file):
// - pcileech_bar_impl_zerowrite4k = zero-initialized read/write BAR.
//     It's possible to modify contents by use of .coe file.
// - pcileech_bar_impl_loopaddr = test core that loops back the 32-bit
//     address of the current read. Does not support writes.
// - pcileech_bar_impl_none = core without any reply.
// 
// (c) Ulf Frisk, 2024
// Author: Ulf Frisk, pcileech@frizk.net
//

`timescale 1ns / 1ps
`include "pcileech_header.svh"

module pcileech_tlps128_bar_controller(
    input                   rst,
    input                   clk,
    input                   bar_en,
    input [15:0]            pcie_id,    
    IfAXIS128.sink_lite     tlps_in,
    IfAXIS128.source        tlps_out,
    output                  int_enable,
    input                   msix_vaild,
    output                  msix_send_done,
    output [31:0]           msix_address,
    output [31:0]           msix_vector,
    input [31:0]            base_address_register,
    input [31:0]            base_address_register_1,
    input [31:0]            base_address_register_2,
    input [31:0]            base_address_register_3,
    input [31:0]            base_address_register_4,
    input [31:0]            base_address_register_5
);
    
    // ------------------------------------------------------------------------
    // 1: TLP RECEIVE:
    // Receive incoming BAR requests from the TLP stream:
    // send them onwards to read and write FIFOs
    // ------------------------------------------------------------------------
    wire in_is_wr_ready;
    bit  in_is_wr_last;
    wire in_is_first    = tlps_in.tuser[0];
    wire in_is_bar      = bar_en && (tlps_in.tuser[8:2] != 0);
    wire in_is_rd       = (in_is_first && tlps_in.tlast && ((tlps_in.tdata[31:25] == 7'b0000000) || (tlps_in.tdata[31:25] == 7'b0010000) || (tlps_in.tdata[31:24] == 8'b00000010)));
    wire in_is_wr       = in_is_wr_last || (in_is_first && in_is_wr_ready && ((tlps_in.tdata[31:25] == 7'b0100000) || (tlps_in.tdata[31:25] == 7'b0110000) || (tlps_in.tdata[31:24] == 8'b01000010)));
    
    always @ ( posedge clk )
        if ( rst ) begin
            in_is_wr_last <= 0;
        end
        else if ( tlps_in.tvalid ) begin
            in_is_wr_last <= !tlps_in.tlast && in_is_wr;
        end

    wire [6:0]  wr_bar;
    wire [31:0] wr_addr;
    wire [3:0]  wr_be;
    wire [31:0] wr_data;
    wire        wr_valid;
    wire [87:0] rd_req_ctx;
    wire [6:0]  rd_req_bar;
    wire [31:0] rd_req_addr;
    wire [3:0]  rd_req_be;
    wire        rd_req_valid;
    wire [87:0] rd_rsp_ctx;
    wire [31:0] rd_rsp_data;
    wire        rd_rsp_valid;
        
    pcileech_tlps128_bar_rdengine i_pcileech_tlps128_bar_rdengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .pcie_id        ( pcie_id                       ),
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_rd ),
        .tlps_out       ( tlps_out                      ),
        // BAR reads:
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_bar     ( rd_req_bar                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_be      ( rd_req_be                     ),
        .rd_req_valid   ( rd_req_valid                  ),
        .rd_rsp_ctx     ( rd_rsp_ctx                    ),
        .rd_rsp_data    ( rd_rsp_data                   ),
        .rd_rsp_valid   ( rd_rsp_valid                  )
    );

    pcileech_tlps128_bar_wrengine i_pcileech_tlps128_bar_wrengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_wr ),
        .tlps_in_ready  ( in_is_wr_ready                ),
        // outgoing BAR writes:
        .wr_bar         ( wr_bar                        ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid                      )
    );
    
    wire [87:0] bar_rsp_ctx[7];
    wire [31:0] bar_rsp_data[7];
    wire        bar_rsp_valid[7];
    
    assign rd_rsp_ctx = bar_rsp_valid[0] ? bar_rsp_ctx[0] :
                        bar_rsp_valid[1] ? bar_rsp_ctx[1] :
                        bar_rsp_valid[2] ? bar_rsp_ctx[2] :
                        bar_rsp_valid[3] ? bar_rsp_ctx[3] :
                        bar_rsp_valid[4] ? bar_rsp_ctx[4] :
                        bar_rsp_valid[5] ? bar_rsp_ctx[5] :
                        bar_rsp_valid[6] ? bar_rsp_ctx[6] : 0;
    assign rd_rsp_data = bar_rsp_valid[0] ? bar_rsp_data[0] :
                        bar_rsp_valid[1] ? bar_rsp_data[1] :
                        bar_rsp_valid[2] ? bar_rsp_data[2] :
                        bar_rsp_valid[3] ? bar_rsp_data[3] :
                        bar_rsp_valid[4] ? bar_rsp_data[4] :
                        bar_rsp_valid[5] ? bar_rsp_data[5] :
                        bar_rsp_valid[6] ? bar_rsp_data[6] : 0;
    assign rd_rsp_valid = bar_rsp_valid[0] || bar_rsp_valid[1] || bar_rsp_valid[2] || bar_rsp_valid[3] || bar_rsp_valid[4] || bar_rsp_valid[5] || bar_rsp_valid[6];
    

    pcileech_bar_impl_zerowrite4k i_bar0(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[0]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[0] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[0]                ),
        .rd_rsp_data    ( bar_rsp_data[0]               ),
        .rd_rsp_valid   ( bar_rsp_valid[0]              )
    );
    
    pcileech_bar_impl_none i_bar1(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[1]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[1] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[1]                ),
        .rd_rsp_data    ( bar_rsp_data[1]               ),
        .rd_rsp_valid   ( bar_rsp_valid[1]              )
    );
    
    pcileech_bar_impl_bar2 i_bar2(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[2]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[2] ),
        .base_address_register( base_address_register_2   ),
        .int_enable     ( int_enable                    ),
        .rd_rsp_ctx     ( bar_rsp_ctx[2]                ),
        .rd_rsp_data    ( bar_rsp_data[2]               ),
        .rd_rsp_valid   ( bar_rsp_valid[2]              )
    );
    
    pcileech_bar_impl_none i_bar3(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[3]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[3] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[3]                ),
        .rd_rsp_data    ( bar_rsp_data[3]               ),
        .rd_rsp_valid   ( bar_rsp_valid[3]              )
    );
    
    pcileech_bar_impl_none i_bar4(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[4]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[4] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[4]                ),
        .rd_rsp_data    ( bar_rsp_data[4]               ),
        .rd_rsp_valid   ( bar_rsp_valid[4]              )
    );
    
    pcileech_bar_impl_none i_bar5(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[5]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[5] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[5]                ),
        .rd_rsp_data    ( bar_rsp_data[5]               ),
        .rd_rsp_valid   ( bar_rsp_valid[5]              )
    );
    
    pcileech_bar_impl_none i_bar6_optrom(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[6]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[6] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[6]                ),
        .rd_rsp_data    ( bar_rsp_data[6]               ),
        .rd_rsp_valid   ( bar_rsp_valid[6]              )
    );


endmodule



// ------------------------------------------------------------------------
// BAR WRITE ENGINE:
// Receives BAR WRITE TLPs and output BAR WRITE requests.
// Holds a 2048-byte buffer.
// Input flow rate is 16bytes/CLK (max).
// Output flow rate is 4bytes/CLK.
// If write engine overflows incoming TLP is completely discarded silently.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_wrengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    output                  tlps_in_ready,
    // outgoing BAR writes:
    output bit [6:0]        wr_bar,
    output bit [31:0]       wr_addr,
    output bit [3:0]        wr_be,
    output bit [31:0]       wr_data,
    output bit              wr_valid
);

    wire            f_rd_en;
    wire [127:0]    f_tdata;
    wire [3:0]      f_tkeepdw;
    wire [8:0]      f_tuser;
    wire            f_tvalid;
    
    bit [127:0]     tdata;
    bit [3:0]       tkeepdw;
    bit             tlast;
    
    bit [3:0]       be_first;
    bit [3:0]       be_last;
    bit             first_dw;
    bit [31:0]      addr;

    fifo_141_141_clk1_bar_wr i_fifo_141_141_clk1_bar_wr(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( {tlps_in.tuser[8:0], tlps_in.tkeepdw, tlps_in.tdata} ),
        .full           (                               ),
        .prog_empty     ( tlps_in_ready                 ),
        .rd_en          ( f_rd_en                       ),
        .dout           ( {f_tuser, f_tkeepdw, f_tdata} ),    
        .empty          (                               ),
        .valid          ( f_tvalid                      )
    );
    
    // STATE MACHINE:
    `define S_ENGINE_IDLE        3'h0
    `define S_ENGINE_FIRST       3'h1
    `define S_ENGINE_4DW_REQDATA 3'h2
    `define S_ENGINE_TX0         3'h4
    `define S_ENGINE_TX1         3'h5
    `define S_ENGINE_TX2         3'h6
    `define S_ENGINE_TX3         3'h7
    (* KEEP = "TRUE" *) bit [3:0] state = `S_ENGINE_IDLE;
    
    assign f_rd_en = (state == `S_ENGINE_IDLE) ||
                     (state == `S_ENGINE_4DW_REQDATA) ||
                     (state == `S_ENGINE_TX3) ||
                     ((state == `S_ENGINE_TX2 && !tkeepdw[3])) ||
                     ((state == `S_ENGINE_TX1 && !tkeepdw[2])) ||
                     ((state == `S_ENGINE_TX0 && !f_tkeepdw[1]));

    always @ ( posedge clk ) begin
        wr_addr     <= addr;
        wr_valid    <= ((state == `S_ENGINE_TX0) && f_tvalid) || (state == `S_ENGINE_TX1) || (state == `S_ENGINE_TX2) || (state == `S_ENGINE_TX3);
        
    end

    always @ ( posedge clk )
        if ( rst ) begin
            state <= `S_ENGINE_IDLE;
        end
        else case ( state )
            `S_ENGINE_IDLE: begin
                state   <= `S_ENGINE_FIRST;
            end
            `S_ENGINE_FIRST: begin
                if ( f_tvalid && f_tuser[0] ) begin
                    wr_bar      <= f_tuser[8:2];
                    tdata       <= f_tdata;
                    tkeepdw     <= f_tkeepdw;
                    tlast       <= f_tuser[1];
                    first_dw    <= 1;
                    be_first    <= f_tdata[35:32];
                    be_last     <= f_tdata[39:36];
                    if ( f_tdata[31:29] == 8'b010 ) begin       // 3 DW header, with data
                        addr    <= { f_tdata[95:66], 2'b00 };
                        state   <= `S_ENGINE_TX3;
                    end
                    else if ( f_tdata[31:29] == 8'b011 ) begin  // 4 DW header, with data
                        addr    <= { f_tdata[127:98], 2'b00 };
                        state   <= `S_ENGINE_4DW_REQDATA;
                    end 
                end
                else begin
                    state   <= `S_ENGINE_IDLE;
                end
            end 
            `S_ENGINE_4DW_REQDATA: begin
                state   <= `S_ENGINE_TX0;
            end
            `S_ENGINE_TX0: begin
                tdata       <= f_tdata;
                tkeepdw     <= f_tkeepdw;
                tlast       <= f_tuser[1];
                addr        <= addr + 4;
                wr_data     <= { f_tdata[0+00+:8], f_tdata[0+08+:8], f_tdata[0+16+:8], f_tdata[0+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (f_tkeepdw[1] ? 4'hf : be_last);
                state       <= f_tvalid ? (f_tkeepdw[1] ? `S_ENGINE_TX1 : `S_ENGINE_FIRST) : `S_ENGINE_IDLE;
            end
            `S_ENGINE_TX1: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[32+00+:8], tdata[32+08+:8], tdata[32+16+:8], tdata[32+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[2] ? 4'hf : be_last);
                state       <= tkeepdw[2] ? `S_ENGINE_TX2 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX2: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[64+00+:8], tdata[64+08+:8], tdata[64+16+:8], tdata[64+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[3] ? 4'hf : be_last);
                state       <= tkeepdw[3] ? `S_ENGINE_TX3 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX3: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[96+00+:8], tdata[96+08+:8], tdata[96+16+:8], tdata[96+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (!tlast ? 4'hf : be_last);
                state       <= !tlast ? `S_ENGINE_TX0 : `S_ENGINE_FIRST;
            end
        endcase

endmodule




// ------------------------------------------------------------------------
// BAR READ ENGINE:
// Receives BAR READ TLPs and output BAR READ requests.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_rdengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    input [15:0]            pcie_id,
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    IfAXIS128.source        tlps_out,
    // BAR reads:
    output [87:0]           rd_req_ctx,
    output [6:0]            rd_req_bar,
    output [31:0]           rd_req_addr,
    output                  rd_req_valid,
    output [3:0]            rd_req_be,        
    input  [87:0]           rd_rsp_ctx,
    input  [31:0]           rd_rsp_data,
    input                   rd_rsp_valid
);
    // ------------------------------------------------------------------------
    // 1: PROCESS AND QUEUE INCOMING READ TLPs:
    // ------------------------------------------------------------------------
    wire [10:0] rd1_in_dwlen    = (tlps_in.tdata[9:0] == 0) ? 11'd1024 : {1'b0, tlps_in.tdata[9:0]};
    wire [6:0]  rd1_in_bar      = tlps_in.tuser[8:2];
    wire [15:0] rd1_in_reqid    = tlps_in.tdata[63:48];
    wire [7:0]  rd1_in_tag      = tlps_in.tdata[47:40];
    wire [31:0] rd1_in_addr     = { ((tlps_in.tdata[31:29] == 3'b000) ? tlps_in.tdata[95:66] : tlps_in.tdata[127:98]), 2'b00 };
    wire [3:0]  rd1_in_be       = tlps_in.tdata[35:32];
    wire [73:0] rd1_in_data;
    assign rd1_in_data[73:63]   = rd1_in_dwlen;
    assign rd1_in_data[62:56]   = rd1_in_bar;   
    assign rd1_in_data[55:48]   = rd1_in_tag;
    assign rd1_in_data[47:32]   = rd1_in_reqid;
    assign rd1_in_data[31:0]    = rd1_in_addr;

    
    wire [3:0]  rd1_out_be;
    wire        rd1_out_be_valid;
    wire        rd1_out_rden;
    wire [73:0] rd1_out_data;
    wire        rd1_out_valid;
    
    fifo_74_74_clk1_bar_rd1 i_fifo_74_74_clk1_bar_rd1(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( rd1_in_data                   ),
        .full           (                               ),
        .rd_en          ( rd1_out_rden                  ),
        .dout           ( rd1_out_data                  ),    
        .empty          (                               ),
        .valid          ( rd1_out_valid                 )
    );
    fifo_4_4_clk1_bar_rd1 i_fifo_4_4_clk1_bar_rd1 (
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( rd1_in_be                     ),
        .full           (                               ),
        .rd_en          ( rd1_out_rden                  ),
        .dout           ( rd1_out_be                    ),
        .empty          (                               ),
        .valid          ( rd1_out_be_valid              )

    );
    
    // ------------------------------------------------------------------------
    // 2: PROCESS AND SPLIT READ TLPs INTO RESPONSE TLP READ REQUESTS AND QUEUE:
    //    (READ REQUESTS LARGER THAN 128-BYTES WILL BE SPLIT INTO MULTIPLE).
    // ------------------------------------------------------------------------
    
    wire [10:0] rd1_out_dwlen       = rd1_out_data[73:63];
    wire [4:0]  rd1_out_dwlen5      = rd1_out_data[67:63];
    wire [4:0]  rd1_out_addr5       = rd1_out_data[6:2];
    
    // 1st "instant" packet:
    wire [4:0]  rd2_pkt1_dwlen_pre  = ((rd1_out_addr5 + rd1_out_dwlen5 > 6'h20) || ((rd1_out_addr5 != 0) && (rd1_out_dwlen5 == 0))) ? (6'h20 - rd1_out_addr5) : rd1_out_dwlen5;
    wire [5:0]  rd2_pkt1_dwlen      = (rd2_pkt1_dwlen_pre == 0) ? 6'h20 : rd2_pkt1_dwlen_pre;
    wire [10:0] rd2_pkt1_dwlen_next = rd1_out_dwlen - rd2_pkt1_dwlen;
    wire        rd2_pkt1_large      = (rd1_out_dwlen > 32) || (rd1_out_dwlen != rd2_pkt1_dwlen);
    wire        rd2_pkt1_tiny       = (rd1_out_dwlen == 1);
    wire [11:0] rd2_pkt1_bc         = rd1_out_dwlen << 2;
    wire [85:0] rd2_pkt1;
    assign      rd2_pkt1[85:74]     = rd2_pkt1_bc;
    assign      rd2_pkt1[73:63]     = rd2_pkt1_dwlen;
    assign      rd2_pkt1[62:0]      = rd1_out_data[62:0];
    
    // Nth packet (if split should take place):
    bit  [10:0] rd2_total_dwlen;
    wire [10:0] rd2_total_dwlen_next = rd2_total_dwlen - 11'h20;
    
    bit  [85:0] rd2_pkt2;
    wire [10:0] rd2_pkt2_dwlen = rd2_pkt2[73:63];
    wire        rd2_pkt2_large = (rd2_total_dwlen > 11'h20);
    
    wire        rd2_out_rden;
    
    // STATE MACHINE:
    `define S2_ENGINE_REQDATA     1'h0
    `define S2_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state2 = `S2_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            state2 <= `S2_ENGINE_REQDATA;
        end
        else case ( state2 )
            `S2_ENGINE_REQDATA: begin
                if ( rd1_out_valid && rd2_pkt1_large ) begin
                    rd2_total_dwlen <= rd2_pkt1_dwlen_next;                             // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_pkt1_dwlen_next << 2;                        // byte-count
                    rd2_pkt2[73:63] <= (rd2_pkt1_dwlen_next > 11'h20) ? 11'h20 : rd2_pkt1_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd1_out_data[62:12];                             // various data
                    rd2_pkt2[11:0]  <= rd1_out_data[11:0] + (rd2_pkt1_dwlen << 2);      // base address (within 4k page)
                    state2 <= `S2_ENGINE_PROCESSING;
                end
            end
            `S2_ENGINE_PROCESSING: begin
                if ( rd2_out_rden ) begin
                    rd2_total_dwlen <= rd2_total_dwlen_next;                                // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_total_dwlen_next << 2;                           // byte-count
                    rd2_pkt2[73:63] <= (rd2_total_dwlen_next > 11'h20) ? 11'h20 : rd2_total_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd2_pkt2[62:12];                                     // various data
                    rd2_pkt2[11:0]  <= rd2_pkt2[11:0] + (rd2_pkt2_dwlen << 2);              // base address (within 4k page)
                    if ( !rd2_pkt2_large ) begin
                        state2 <= `S2_ENGINE_REQDATA;
                    end
                end
            end
        endcase
    
    assign rd1_out_rden = rd2_out_rden && (((state2 == `S2_ENGINE_REQDATA) && (!rd1_out_valid || rd2_pkt1_tiny)) || ((state2 == `S2_ENGINE_PROCESSING) && !rd2_pkt2_large));

    wire [85:0] rd2_in_data  = (state2 == `S2_ENGINE_REQDATA) ? rd2_pkt1 : rd2_pkt2;
    wire        rd2_in_valid = rd1_out_valid || ((state2 == `S2_ENGINE_PROCESSING) && rd2_out_rden);
    wire [3:0]  rd2_in_be       = rd1_out_be;
    wire        rd2_in_be_valid = rd1_out_valid;

    bit  [85:0] rd2_out_data;
    bit         rd2_out_valid;
    bit  [3:0]  rd2_out_be;
    bit         rd2_out_be_valid;
    always @ ( posedge clk ) begin
        rd2_out_data    <= rd2_in_valid ? rd2_in_data : rd2_out_data;
        rd2_out_valid   <= rd2_in_valid && !rst;
        rd2_out_be       <= rd2_in_be_valid ? rd2_in_be : rd2_out_data;
        rd2_out_be_valid <= rd2_in_be_valid && !rst;  
    end

    // ------------------------------------------------------------------------
    // 3: PROCESS EACH READ REQUEST PACKAGE PER INDIVIDUAL 32-bit READ DWORDS:
    // ------------------------------------------------------------------------

    wire [4:0]  rd2_out_dwlen   = rd2_out_data[67:63];
    wire        rd2_out_last    = (rd2_out_dwlen == 1);
    wire [9:0]  rd2_out_dwaddr  = rd2_out_data[11:2];
    
    wire        rd3_enable;
    
    bit [3:0]   rd3_process_be;
    bit         rd3_process_valid;
    bit         rd3_process_first;
    bit         rd3_process_last;
    bit [4:0]   rd3_process_dwlen;
    bit [9:0]   rd3_process_dwaddr;
    bit [85:0]  rd3_process_data;
    wire        rd3_process_next_last = (rd3_process_dwlen == 2);
    wire        rd3_process_nextnext_last = (rd3_process_dwlen <= 3);
    assign rd_req_be    = rd3_process_be;
    assign rd_req_ctx   = { rd3_process_first, rd3_process_last, rd3_process_data };
    assign rd_req_bar   = rd3_process_data[62:56];
    assign rd_req_addr  = { rd3_process_data[31:12], rd3_process_dwaddr, 2'b00 };
    assign rd_req_valid = rd3_process_valid;
    
    // STATE MACHINE:
    `define S3_ENGINE_REQDATA     1'h0
    `define S3_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state3 = `S3_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            rd3_process_valid   <= 1'b0;
            state3              <= `S3_ENGINE_REQDATA;
        end
        else case ( state3 )
            `S3_ENGINE_REQDATA: begin
                if ( rd2_out_valid ) begin
                    rd3_process_valid       <= 1'b1;
                    rd3_process_first       <= 1'b1;                    // FIRST
                    rd3_process_last        <= rd2_out_last;            // LAST (low 5 bits of dwlen == 1, [max pktlen = 0x20))
                    rd3_process_dwlen       <= rd2_out_dwlen;           // PKT LENGTH IN DW
                    rd3_process_dwaddr      <= rd2_out_dwaddr;          // DWADDR OF THIS DWORD
                    rd3_process_data[85:0]  <= rd2_out_data[85:0];      // FORWARD / SAVE DATA
                    if ( rd2_out_be_valid ) begin
                        rd3_process_be <= rd2_out_be;
                    end else begin
                        rd3_process_be <= 4'hf;
                    end
                    if ( !rd2_out_last ) begin
                        state3 <= `S3_ENGINE_PROCESSING;
                    end
                end
                else begin
                    rd3_process_valid       <= 1'b0;
                end
            end
            `S3_ENGINE_PROCESSING: begin
                rd3_process_first           <= 1'b0;                    // FIRST
                rd3_process_last            <= rd3_process_next_last;   // LAST
                rd3_process_dwlen           <= rd3_process_dwlen - 1;   // LEN DEC
                rd3_process_dwaddr          <= rd3_process_dwaddr + 1;  // ADDR INC
                if ( rd3_process_next_last ) begin
                    state3 <= `S3_ENGINE_REQDATA;
                end
            end
        endcase

    assign rd2_out_rden = rd3_enable && (
        ((state3 == `S3_ENGINE_REQDATA) && (!rd2_out_valid || rd2_out_last)) ||
        ((state3 == `S3_ENGINE_PROCESSING) && rd3_process_nextnext_last));
    
    // ------------------------------------------------------------------------
    // 4: PROCESS RESPONSES:
    // ------------------------------------------------------------------------
    
    wire        rd_rsp_first    = rd_rsp_ctx[87];
    wire        rd_rsp_last     = rd_rsp_ctx[86];
    
    wire [9:0]  rd_rsp_dwlen    = rd_rsp_ctx[72:63];
    wire [11:0] rd_rsp_bc       = rd_rsp_ctx[85:74];
    wire [15:0] rd_rsp_reqid    = rd_rsp_ctx[47:32];
    wire [7:0]  rd_rsp_tag      = rd_rsp_ctx[55:48];
    wire [6:0]  rd_rsp_lowaddr  = rd_rsp_ctx[6:0];
    wire [31:0] rd_rsp_addr     = rd_rsp_ctx[31:0];
    wire [31:0] rd_rsp_data_bs  = { rd_rsp_data[7:0], rd_rsp_data[15:8], rd_rsp_data[23:16], rd_rsp_data[31:24] };
    
    // 1: 32-bit -> 128-bit state machine:
    bit [127:0] tdata;
    bit [3:0]   tkeepdw = 0;
    bit         tlast;
    bit         first   = 1;
    wire        tvalid  = tlast || tkeepdw[3];
    
    always @ ( posedge clk )
        if ( rst ) begin
            tkeepdw <= 0;
            tlast   <= 0;
            first   <= 0;
        end
        else if ( rd_rsp_valid && rd_rsp_first ) begin
            tkeepdw         <= 4'b1111;
            tlast           <= rd_rsp_last;
            first           <= 1'b1;
            tdata[31:0]     <= { 22'b0100101000000000000000, rd_rsp_dwlen };            // format, type, length
            tdata[63:32]    <= { pcie_id[7:0], pcie_id[15:8], 4'b0, rd_rsp_bc };        // pcie_id, byte_count
            tdata[95:64]    <= { rd_rsp_reqid, rd_rsp_tag, 1'b0, rd_rsp_lowaddr };      // req_id, tag, lower_addr
            tdata[127:96]   <= rd_rsp_data_bs;
        end
        else begin
            tlast   <= rd_rsp_valid && rd_rsp_last;
            tkeepdw <= tvalid ? (rd_rsp_valid ? 4'b0001 : 4'b0000) : (rd_rsp_valid ? ((tkeepdw << 1) | 1'b1) : tkeepdw);
            first   <= 0;
            if ( rd_rsp_valid ) begin
                if ( tvalid || !tkeepdw[0] )
                    tdata[31:0]   <= rd_rsp_data_bs;
                if ( !tkeepdw[1] )
                    tdata[63:32]  <= rd_rsp_data_bs;
                if ( !tkeepdw[2] )
                    tdata[95:64]  <= rd_rsp_data_bs;
                if ( !tkeepdw[3] )
                    tdata[127:96] <= rd_rsp_data_bs;   
            end
        end
    
    // 2.1 - submit to output fifo - will feed into mux/pcie core.
    fifo_134_134_clk1_bar_rdrsp i_fifo_134_134_clk1_bar_rdrsp(
        .srst           ( rst                       ),
        .clk            ( clk                       ),
        .din            ( { first, tlast, tkeepdw, tdata } ),
        .wr_en          ( tvalid                    ),
        .rd_en          ( tlps_out.tready           ),
        .dout           ( { tlps_out.tuser[0], tlps_out.tlast, tlps_out.tkeepdw, tlps_out.tdata } ),
        .full           (                           ),
        .empty          (                           ),
        .prog_empty     ( rd3_enable                ),
        .valid          ( tlps_out.tvalid           )
    );
    
    assign tlps_out.tuser[1] = tlps_out.tlast;
    assign tlps_out.tuser[8:2] = 0;
    
    // 2.2 - packet count:
    bit [10:0]  pkt_count       = 0;
    wire        pkt_count_dec   = tlps_out.tvalid && tlps_out.tlast;
    wire        pkt_count_inc   = tvalid && tlast;
    wire [10:0] pkt_count_next  = pkt_count + pkt_count_inc - pkt_count_dec;
    assign tlps_out.has_data    = (pkt_count_next > 0);
    
    always @ ( posedge clk ) begin
        pkt_count <= rst ? 0 : pkt_count_next;
    end

endmodule


// ------------------------------------------------------------------------
// Example BAR implementation that does nothing but drop any read/writes
// silently without generating a response.
// This is only recommended for placeholder designs.
// Latency = N/A.
// ------------------------------------------------------------------------
module pcileech_bar_impl_none(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    initial rd_rsp_ctx = 0;
    initial rd_rsp_data = 0;
    initial rd_rsp_valid = 0;

endmodule




// ------------------------------------------------------------------------
// Example BAR implementation of "address loopback" which can be useful
// for testing. Any read to a specific BAR address will result in the
// address as response.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_loopaddr(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input [87:0]        rd_req_ctx,
    input [31:0]        rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]      rd_req_ctx_1;
    bit [31:0]      rd_req_addr_1;
    bit             rd_req_valid_1;
    
    always @ ( posedge clk ) begin
        rd_req_ctx_1    <= rd_req_ctx;
        rd_req_addr_1   <= rd_req_addr;
        rd_req_valid_1  <= rd_req_valid;
        rd_rsp_ctx      <= rd_req_ctx_1;
        rd_rsp_data     <= rd_req_addr_1;
        rd_rsp_valid    <= rd_req_valid_1;
    end    

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of a 4kB writable initial-zero BAR.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_zerowrite4k(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]  drd_req_ctx;
    bit         drd_req_valid;
    wire [31:0] doutb;
    
    always @ ( posedge clk ) begin
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        rd_rsp_data     <= doutb; 
    end
    
    bram_bar_zero4k i_bram_bar_zero4k(
        // Port A - write:
        .addra  ( wr_addr[11:2]     ),
        .clka   ( clk               ),
        .dina   ( wr_data           ),
        .ena    ( wr_valid          ),
        .wea    ( wr_be             ),
        // Port A - read (2 CLK latency):
        .addrb  ( rd_req_addr[11:2] ),
        .clkb   ( clk               ),
        .doutb  ( doutb             ),
        .enb    ( rd_req_valid      )
    );

endmodule


`define MAC_RANDOM_NUM1 13
`define MAC_RANDOM_NUM2 2
`define MAC_RANDOM_NUM3 13
`define MAC_RANDOM_NUM4 9
`define MAC_RANDOM_NUM5 7
`define MAC_RANDOM_NUM6 5


module pcileech_bar_impl_bar2(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    input  [31:0]       base_address_register,
    // outgoing BAR read replies:
    output wire         int_enable,
    output reg [87:0]   rd_rsp_ctx,
    output reg [31:0]   rd_rsp_data,
    output reg          rd_rsp_valid
);
                     
    reg [87:0]      drd_req_ctx;
    reg [31:0]      drd_req_addr;
    reg             drd_req_valid;
                  
    reg [31:0]      dwr_addr;
    reg [31:0]      dwr_data;
    reg             dwr_valid;
               
    reg [31:0]      data_32;
              
    time number = 0;

    assign int_enable = 1'b1;
                  
    always @ (posedge clk) begin
        if (rst)
            number <= 0;
               
        number          <= number + 1;
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        dwr_valid       <= wr_valid;
        drd_req_addr    <= rd_req_addr;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        dwr_addr        <= wr_addr;
        dwr_data        <= wr_data;

        if (drd_req_valid) begin
            case (({drd_req_addr[31:24], drd_req_addr[23:16], drd_req_addr[15:08], drd_req_addr[07:00]} - (base_address_register & 32'hFFFFFFF0)) & 32'hFFFF)
                16'h0000 : rd_rsp_data <= 32'hFDC3B2D2;
                16'h0004 : rd_rsp_data <= 32'h15030012;
                16'h0008 : rd_rsp_data <= 32'h00207C2B;
                16'h0010 : rd_rsp_data <= 32'h4007EB03;
                16'h0014 : rd_rsp_data <= 32'h10562175;
                16'h0018 : rd_rsp_data <= 32'h00400100;
                16'h001C : rd_rsp_data <= 32'h07F6E100;
                16'h0020 : rd_rsp_data <= 32'h05010101;
                16'h0024 : rd_rsp_data <= 32'h000F81F9;
                16'h0028 : rd_rsp_data <= 32'hF4004783;
                16'h002C : rd_rsp_data <= 32'hF0AAA596;
                16'h0030 : rd_rsp_data <= 32'hF261FAFF;
                16'h0034 : rd_rsp_data <= 32'h34000000;
                16'h0040 : rd_rsp_data <= 32'h00000220;
                16'h0044 : rd_rsp_data <= 32'h00200090;
                16'h0048 : rd_rsp_data <= 32'h00020000;
                16'h004C : rd_rsp_data <= 32'h0FE28282;
                16'h0050 : rd_rsp_data <= 32'h80000000;
                16'h0060 : rd_rsp_data <= 32'h00000062;
                16'h0064 : rd_rsp_data <= 32'h30030104;
                16'h0068 : rd_rsp_data <= 32'h80086804;
                16'h006C : rd_rsp_data <= 32'h000000E0;
                16'h0074 : rd_rsp_data <= 32'h00000405;
                16'h0078 : rd_rsp_data <= 32'h0A1E002A;
                16'h007C : rd_rsp_data <= 32'h00000083;
                16'h0080 : rd_rsp_data <= 32'h800706C6;
                16'h0090 : rd_rsp_data <= 32'hD5000000;
                16'h0094 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00A0 : rd_rsp_data <= 32'h00000620;
                16'h00A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00A8 : rd_rsp_data <= 32'hFF000000;
                16'h00AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00B0 : rd_rsp_data <= 32'h31000603;
                16'h00B4 : rd_rsp_data <= 32'h00100041;
                16'h00B8 : rd_rsp_data <= 32'h10000F00;
                16'h00C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00CC : rd_rsp_data <= 32'h00000029;
                16'h00D0 : rd_rsp_data <= 32'h001FC002;
                16'h00DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h00F0 : rd_rsp_data <= 32'h0C44113B;
                16'h00F4 : rd_rsp_data <= 32'h0000006B;
                16'h00F8 : rd_rsp_data <= 32'h00038129;
                16'h00FC : rd_rsp_data <= 32'h00000207;
                16'h0100 : rd_rsp_data <= 32'h000006FF;
                16'h0104 : rd_rsp_data <= 32'h00000020;
                16'h010C : rd_rsp_data <= 32'h0000F5B1;
                16'h0114 : rd_rsp_data <= 32'h3CFF0FF5;
                16'h011C : rd_rsp_data <= 32'h11981198;
                16'h0130 : rd_rsp_data <= 32'h72070012;
                16'h0134 : rd_rsp_data <= 32'h00000009;
                16'h0138 : rd_rsp_data <= 32'hE213091F;
                16'h013C : rd_rsp_data <= 32'h10000200;
                16'h0164 : rd_rsp_data <= 32'h00000001;
                16'h0174 : rd_rsp_data <= 32'h000008FF;
                16'h0194 : rd_rsp_data <= 32'h10000001;
                16'h0198 : rd_rsp_data <= 32'h000B0047;
                16'h01C4 : rd_rsp_data <= 32'hFE0057FC;
                16'h01D0 : rd_rsp_data <= 32'h00FF0F1E;
                16'h01D4 : rd_rsp_data <= 32'h00FF0F1E;
                16'h01D8 : rd_rsp_data <= 32'h00FF001E;
                16'h01DC : rd_rsp_data <= 32'h00FF001E;
                16'h01E4 : rd_rsp_data <= 32'h00000523;
                16'h01E8 : rd_rsp_data <= 32'h00000880;
                16'h01EC : rd_rsp_data <= 32'hB0000C1C;
                16'h0200 : rd_rsp_data <= 32'h00E40808;
                16'h0204 : rd_rsp_data <= 32'h00E40808;
                16'h0208 : rd_rsp_data <= 32'h6B00F510;
                16'h020C : rd_rsp_data <= 32'h00FD0000;
                16'h0224 : rd_rsp_data <= 32'h00002020;
                16'h0228 : rd_rsp_data <= 32'h0000F500;
                16'h0280 : rd_rsp_data <= 32'h00002003;
                16'h0284 : rd_rsp_data <= 32'h00020000;
                16'h0290 : rd_rsp_data <= 32'h00000004;
                16'h0294 : rd_rsp_data <= 32'h00003D00;
                16'h0300 : rd_rsp_data <= 32'hA7038000;
                16'h0308 : rd_rsp_data <= 32'h7013C000;
                16'h0310 : rd_rsp_data <= 32'h70069000;
                16'h0318 : rd_rsp_data <= 32'h700CB000;
                16'h0320 : rd_rsp_data <= 32'h700DD000;
                16'h0328 : rd_rsp_data <= 32'h700FC000;
                16'h0330 : rd_rsp_data <= 32'h70146000;
                16'h0338 : rd_rsp_data <= 32'h6E9C7000;
                16'h0340 : rd_rsp_data <= 32'h70050000;
                16'h0380 : rd_rsp_data <= 32'hA2001200;
                16'h0384 : rd_rsp_data <= 32'h12001200;
                16'h0388 : rd_rsp_data <= 32'h12001200;
                16'h038C : rd_rsp_data <= 32'h12001200;
                16'h0390 : rd_rsp_data <= 32'h12001200;
                16'h0394 : rd_rsp_data <= 32'h12001200;
                16'h0398 : rd_rsp_data <= 32'h12001200;
                16'h039C : rd_rsp_data <= 32'h401D401D;
                16'h03B0 : rd_rsp_data <= 32'h01600160;
                16'h03B4 : rd_rsp_data <= 32'h00730073;
                16'h03D8 : rd_rsp_data <= 32'h08008004;
                16'h03E8 : rd_rsp_data <= 32'h97020D00;
                16'h03EC : rd_rsp_data <= 32'h00020D00;
                16'h03F0 : rd_rsp_data <= 32'h04000718;
                16'h03F4 : rd_rsp_data <= 32'h6FB76FB7;
                16'h03F8 : rd_rsp_data <= 32'h0000000A;
                16'h0400 : rd_rsp_data <= 32'h007F80FF;
                16'h0404 : rd_rsp_data <= 32'h007F80FF;
                16'h0408 : rd_rsp_data <= 32'h007F80FF;
                16'h040C : rd_rsp_data <= 32'h007F80FF;
                16'h0410 : rd_rsp_data <= 32'h027F80FF;
                16'h0414 : rd_rsp_data <= 32'h007F80FF;
                16'h0418 : rd_rsp_data <= 32'h0FFF00F5;
                16'h041C : rd_rsp_data <= 32'h000000F5;
                16'h0420 : rd_rsp_data <= 32'hFF711F80;
                16'h0424 : rd_rsp_data <= 32'h6A30F5F5;
                16'h0428 : rd_rsp_data <= 32'h07070E10;
                16'h0430 : rd_rsp_data <= 32'h01000000;
                16'h0434 : rd_rsp_data <= 32'h07060504;
                16'h0438 : rd_rsp_data <= 32'h01000000;
                16'h043C : rd_rsp_data <= 32'h07060504;
                16'h0440 : rd_rsp_data <= 32'h00000FFF;
                16'h0444 : rd_rsp_data <= 32'h00000010;
                16'h0448 : rd_rsp_data <= 32'h3E0FF000;
                16'h044C : rd_rsp_data <= 32'h00000010;
                16'h0450 : rd_rsp_data <= 32'h000FF000;
                16'h0454 : rd_rsp_data <= 32'hF55E0000;
                16'h0458 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h045C : rd_rsp_data <= 32'h1000F500;
                16'h0460 : rd_rsp_data <= 32'h03086666;
                16'h0464 : rd_rsp_data <= 32'h00FF00FF;
                16'h0468 : rd_rsp_data <= 32'h007F80FF;
                16'h046C : rd_rsp_data <= 32'h007F80FF;
                16'h0470 : rd_rsp_data <= 32'h007F80FF;
                16'h0474 : rd_rsp_data <= 32'h007F80FF;
                16'h0480 : rd_rsp_data <= 32'h000C0400;
                16'h04AC : rd_rsp_data <= 32'h12010200;
                16'h04B0 : rd_rsp_data <= 32'h40404040;
                16'h04BC : rd_rsp_data <= 32'h00040040;
                16'h04C0 : rd_rsp_data <= 32'h10001000;
                16'h04C4 : rd_rsp_data <= 32'h80040340;
                16'h04C8 : rd_rsp_data <= 32'h171708FF;
                16'h04CC : rd_rsp_data <= 32'h0201FF7F;
                16'h04DC : rd_rsp_data <= 32'h00000160;
                16'h04E4 : rd_rsp_data <= 32'h25240C0C;
                16'h04E8 : rd_rsp_data <= 32'h06060606;
                16'h04F0 : rd_rsp_data <= 32'h0000C100;
                16'h04F4 : rd_rsp_data <= 32'h00200001;
                16'h04FC : rd_rsp_data <= 32'hFFFF0000;
                16'h0500 : rd_rsp_data <= 32'h002F3210;
                16'h0504 : rd_rsp_data <= 32'h0000A422;
                16'h0508 : rd_rsp_data <= 32'h005EA42B;
                16'h050C : rd_rsp_data <= 32'h0000A422;
                16'h0510 : rd_rsp_data <= 32'h28004413;
                16'h0514 : rd_rsp_data <= 32'h0E100E10;
                16'h0518 : rd_rsp_data <= 32'h0916FE00;
                16'h0520 : rd_rsp_data <= 32'h00003F0F;
                16'h0524 : rd_rsp_data <= 32'h21FF4F0F;
                16'h0528 : rd_rsp_data <= 32'h806C0A8F;
                16'h0540 : rd_rsp_data <= 32'h8000FF12;
                16'h0544 : rd_rsp_data <= 32'h00400180;
                16'h0550 : rd_rsp_data <= 32'h0000001D;
                16'h0554 : rd_rsp_data <= 32'h00640064;
                16'h0558 : rd_rsp_data <= 32'h00020202;
                16'h055C : rd_rsp_data <= 32'h0F0FFF50;
                16'h0560 : rd_rsp_data <= 32'h0C4020FA;
                16'h0568 : rd_rsp_data <= 32'h0C402109;
                16'h0570 : rd_rsp_data <= 32'h000A0002;
                16'h0574 : rd_rsp_data <= 32'h03FF1000;
                16'h058C : rd_rsp_data <= 32'h06200060;
                16'h0590 : rd_rsp_data <= 32'h000F000F;
                16'h05A0 : rd_rsp_data <= 32'h02020202;
                16'h05A4 : rd_rsp_data <= 32'h00010202;
                16'h05CC : rd_rsp_data <= 32'h11E21051;
                16'h05E0 : rd_rsp_data <= 32'h00001000;
                16'h05E4 : rd_rsp_data <= 32'h00003000;
                16'h05E8 : rd_rsp_data <= 32'h00001000;
                16'h05EC : rd_rsp_data <= 32'h00000003;
                16'h05FC : rd_rsp_data <= 32'hFFFF0000;
                16'h0600 : rd_rsp_data <= 32'h04000000;
                16'h0604 : rd_rsp_data <= 32'h00003000;
                16'h0608 : rd_rsp_data <= 32'hF000780E;
                16'h060C : rd_rsp_data <= 32'h04000420;
                // 这里是模拟了一个随机MAC 但是这只是寄存器映射 实际网卡的MAC是从Efuse取出 所以这里是无效的
//                16'h0610 : begin
//                        rd_rsp_data[7:0]   <= 8'h00;
//                        rd_rsp_data[15:8]  <= 8'h0C;
//                        rd_rsp_data[23:16] <= 8'h43;
//                        rd_rsp_data[31:24] <= ((0 + (number + `MAC_RANDOM_NUM1) % (15 + 1 - 0)) << 4) | (0 + (number + `MAC_RANDOM_NUM2) % (15 + 1 - 0)); 
//                end
//                16'h0614 : begin
//                        rd_rsp_data[7:0]   <= ((0 + (number + `MAC_RANDOM_NUM3) % (15 + 1 - 0)) << 4) | (0 + (number + `MAC_RANDOM_NUM6) % (15 + 1 - 0));
//                        rd_rsp_data[15:8]  <= ((0 + (number + `MAC_RANDOM_NUM5) % (15 + 1 - 0)) << 4) | (0 + (number + `MAC_RANDOM_NUM6) % (15 + 1 - 0));
//                        rd_rsp_data[31:16] <= 16'h0000;
//                end
                16'h0610 : rd_rsp_data <= 32'h04430C00;
                16'h0614 : rd_rsp_data <= 32'h0000EB39;
                16'h0620 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0624 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0638 : rd_rsp_data <= 32'h0E102850;
                16'h063C : rd_rsp_data <= 32'h0E0E0A0A;
                16'h0640 : rd_rsp_data <= 32'h00401440;
                16'h0650 : rd_rsp_data <= 32'h00EB0426;
                16'h0658 : rd_rsp_data <= 32'hFFFFFFFF;
                16'h065C : rd_rsp_data <= 32'hFFFFFFFF;
                16'h0660 : rd_rsp_data <= 32'h00810010;
                16'h0664 : rd_rsp_data <= 32'h00000005;
                16'h0668 : rd_rsp_data <= 32'h0E301000;
                16'h066C : rd_rsp_data <= 32'h00052000;
                16'h0670 : rd_rsp_data <= 32'h000100FF;
                16'h0680 : rd_rsp_data <= 32'h000000EC;
                16'h0690 : rd_rsp_data <= 32'h000F0000;
                16'h0694 : rd_rsp_data <= 32'h000A0200;
                16'h06A4 : rd_rsp_data <= 32'h0000FFFF;
                16'h06B8 : rd_rsp_data <= 32'h00000008;
                16'h06D8 : rd_rsp_data <= 32'h0000003F;
                16'h0700 : rd_rsp_data <= 32'h04430C02;
                16'h0704 : rd_rsp_data <= 32'h0000EB39;
                16'h0708 : rd_rsp_data <= 32'h87654321;
                16'h0718 : rd_rsp_data <= 32'h20000200;
                16'h0750 : rd_rsp_data <= 32'h00000076;
                16'h0778 : rd_rsp_data <= 32'h00000001;
                16'h0794 : rd_rsp_data <= 32'h0000017F;
                16'h0798 : rd_rsp_data <= 32'h88E088E0;
                16'h079C : rd_rsp_data <= 32'h880B880B;
                16'h07A0 : rd_rsp_data <= 32'h06492A30;
                16'h07A4 : rd_rsp_data <= 32'h0B6F27C2;
                16'h07A8 : rd_rsp_data <= 32'h804040AA;
                16'h0800 : rd_rsp_data <= 32'h83040000;
                16'h0804 : rd_rsp_data <= 32'h00000003;
                16'h0808 : rd_rsp_data <= 32'h0000FC00;
                16'h080C : rd_rsp_data <= 32'h0000000A;
                16'h0810 : rd_rsp_data <= 32'h10001331;
                16'h0814 : rd_rsp_data <= 32'h020C3D10;
                16'h0818 : rd_rsp_data <= 32'h02220385;
                16'h0820 : rd_rsp_data <= 32'h01000100;
                16'h0824 : rd_rsp_data <= 32'hA1390204;
                16'h0828 : rd_rsp_data <= 32'h01000100;
                16'h082C : rd_rsp_data <= 32'h0C390204;
                16'h0830 : rd_rsp_data <= 32'h29292929;
                16'h0834 : rd_rsp_data <= 32'h29292929;
                16'h0838 : rd_rsp_data <= 32'h23232330;
                16'h083C : rd_rsp_data <= 32'h2B2B2B2B;
                16'h0840 : rd_rsp_data <= 32'h04237CE8;
                16'h0844 : rd_rsp_data <= 32'h01807C0A;
                16'h0848 : rd_rsp_data <= 32'h292B2B2B;
                16'h084C : rd_rsp_data <= 32'h29292929;
                16'h0858 : rd_rsp_data <= 32'h009A009A;
                16'h085C : rd_rsp_data <= 32'h01000014;
                16'h0860 : rd_rsp_data <= 32'h66F60010;
                16'h0864 : rd_rsp_data <= 32'h061F0010;
                16'h0868 : rd_rsp_data <= 32'h27292929;
                16'h086C : rd_rsp_data <= 32'h23232323;
                16'h0874 : rd_rsp_data <= 32'h55004200;
                16'h0878 : rd_rsp_data <= 32'h08080808;
                16'h0880 : rd_rsp_data <= 32'hB0000C1C;
                16'h0884 : rd_rsp_data <= 32'h00000001;
                16'h088C : rd_rsp_data <= 32'hCC0000C0;
                16'h0890 : rd_rsp_data <= 32'h605C0903;
                16'h0894 : rd_rsp_data <= 32'hFFFEFFFF;
                16'h0898 : rd_rsp_data <= 32'h44403C38;
                16'h089C : rd_rsp_data <= 32'h54504C48;
                16'h08A0 : rd_rsp_data <= 32'h00100000;
                16'h08A4 : rd_rsp_data <= 32'h00100000;
                16'h08A8 : rd_rsp_data <= 32'h0000010F;
                16'h08AC : rd_rsp_data <= 32'h00001C80;
                16'h08B4 : rd_rsp_data <= 32'h00030000;
                16'h08B8 : rd_rsp_data <= 32'h00107CE8;
                16'h08BC : rd_rsp_data <= 32'h00107C0A;
                16'h08C4 : rd_rsp_data <= 32'h00000B82;
                16'h08D0 : rd_rsp_data <= 32'h0000342D;
                16'h08D4 : rd_rsp_data <= 32'h0000CBD4;
                16'h08D8 : rd_rsp_data <= 32'h04010100;
                16'h08DC : rd_rsp_data <= 32'h01146E3F;
                16'h08E0 : rd_rsp_data <= 32'h02040204;
                16'h08E8 : rd_rsp_data <= 32'hF802070C;
                16'h08EC : rd_rsp_data <= 32'h29292929;
                16'h08F0 : rd_rsp_data <= 32'h29292929;
                16'h08F4 : rd_rsp_data <= 32'h80000000;
                16'h08F8 : rd_rsp_data <= 32'h00001818;
                16'h0904 : rd_rsp_data <= 32'h00000023;
                16'h0908 : rd_rsp_data <= 32'h00000208;
                16'h090C : rd_rsp_data <= 32'h81121313;
                16'h0910 : rd_rsp_data <= 32'h806C0001;
                16'h0914 : rd_rsp_data <= 32'h00000001;
                16'h091C : rd_rsp_data <= 32'h00010000;
                16'h0924 : rd_rsp_data <= 32'h00000001;
                16'h094C : rd_rsp_data <= 32'h00000008;
                16'h09C0 : rd_rsp_data <= 32'h002A513E;
                16'h09C4 : rd_rsp_data <= 32'h005B3FF5;
                16'h0A00 : rd_rsp_data <= 32'h00D047C8;
                16'h0A04 : rd_rsp_data <= 32'h81FF800C;
                16'h0A08 : rd_rsp_data <= 32'h9C408300;
                16'h0A0C : rd_rsp_data <= 32'h2E68120F;
                16'h0A10 : rd_rsp_data <= 32'h95009B78;
                16'h0A14 : rd_rsp_data <= 32'h1114D028;
                16'h0A18 : rd_rsp_data <= 32'h00881117;
                16'h0A1C : rd_rsp_data <= 32'h89140F00;
                16'h0A20 : rd_rsp_data <= 32'h1A1B0010;
                16'h0A24 : rd_rsp_data <= 32'h090E1317;
                16'h0A28 : rd_rsp_data <= 32'h00000204;
                16'h0A2C : rd_rsp_data <= 32'h00D3A000;
                16'h0A30 : rd_rsp_data <= 32'h00000001;
                16'h0A38 : rd_rsp_data <= 32'h00000001;
                16'h0A3C : rd_rsp_data <= 32'h00000006;
                16'h0A40 : rd_rsp_data <= 32'h000000F8;
                16'h0A44 : rd_rsp_data <= 32'h000000F6;
                16'h0A48 : rd_rsp_data <= 32'h00000009;
                16'h0A50 : rd_rsp_data <= 32'h630FE880;
                16'h0A54 : rd_rsp_data <= 32'h8030B3FC;
                16'h0A58 : rd_rsp_data <= 32'h02005881;
                16'h0A5C : rd_rsp_data <= 32'h0000043F;
                16'h0A60 : rd_rsp_data <= 32'h8080A903;
                16'h0A70 : rd_rsp_data <= 32'h101FFF00;
                16'h0A74 : rd_rsp_data <= 32'h00000007;
                16'h0A78 : rd_rsp_data <= 32'h00000900;
                16'h0A7C : rd_rsp_data <= 32'h225B0606;
                16'h0A80 : rd_rsp_data <= 32'h218075B1;
                16'h0AB0 : rd_rsp_data <= 32'h000000F9;
                16'h0B68 : rd_rsp_data <= 32'h80000000;
                16'h0B6C : rd_rsp_data <= 32'h80000000;
                16'h0BD8 : rd_rsp_data <= 32'h0283000F;
                16'h0BDC : rd_rsp_data <= 32'h01000000;
                16'h0BE0 : rd_rsp_data <= 32'h01000000;
                16'h0BE4 : rd_rsp_data <= 32'h01000000;
                16'h0BE8 : rd_rsp_data <= 32'h01000000;
                16'h0BEC : rd_rsp_data <= 32'h01000000;
                16'h0BF0 : rd_rsp_data <= 32'h01000000;
                16'h0BF4 : rd_rsp_data <= 32'h01000000;
                16'h0BF8 : rd_rsp_data <= 32'h01000000;
                16'h0C00 : rd_rsp_data <= 32'h48071D40;
                16'h0C04 : rd_rsp_data <= 32'h03A05633;
                16'h0C08 : rd_rsp_data <= 32'h000000E4;
                16'h0C0C : rd_rsp_data <= 32'h6C6C6C6C;
                16'h0C10 : rd_rsp_data <= 32'h08800000;
                16'h0C14 : rd_rsp_data <= 32'h4000E907;
                16'h0C18 : rd_rsp_data <= 32'h08800000;
                16'h0C1C : rd_rsp_data <= 32'h40000105;
                16'h0C30 : rd_rsp_data <= 32'h69E9AC47;
                16'h0C34 : rd_rsp_data <= 32'h469652AF;
                16'h0C38 : rd_rsp_data <= 32'h49795994;
                16'h0C3C : rd_rsp_data <= 32'h0A97971C;
                16'h0C40 : rd_rsp_data <= 32'h1F7C403F;
                16'h0C44 : rd_rsp_data <= 32'h000100B7;
                16'h0C48 : rd_rsp_data <= 32'hEC020107;
                16'h0C4C : rd_rsp_data <= 32'h00F603FD;
                16'h0C50 : rd_rsp_data <= 32'h0004002A;
                16'h0C54 : rd_rsp_data <= 32'h0080801F;
                16'h0C58 : rd_rsp_data <= 32'h0000002A;
                16'h0C5C : rd_rsp_data <= 32'h00248492;
                16'h0C64 : rd_rsp_data <= 32'h2112848B;
                16'h0C68 : rd_rsp_data <= 32'h47C00BFF;
                16'h0C6C : rd_rsp_data <= 32'h00000036;
                16'h0C70 : rd_rsp_data <= 32'h00000600;
                16'h0C74 : rd_rsp_data <= 32'h02013269;
                16'h0C78 : rd_rsp_data <= 32'h407F0001;
                16'h0C7C : rd_rsp_data <= 32'h00B91612;
                16'h0C80 : rd_rsp_data <= 32'h400100FE;
                16'h0C84 : rd_rsp_data <= 32'h21F60000;
                16'h0C88 : rd_rsp_data <= 32'h40040100;
                16'h0C8C : rd_rsp_data <= 32'hA0E40000;
                16'h0C90 : rd_rsp_data <= 32'h00121820;
                16'h0C98 : rd_rsp_data <= 32'h00121820;
                16'h0C9C : rd_rsp_data <= 32'h00007F7F;
                16'h0CA0 : rd_rsp_data <= 32'hF0000000;
                16'h0CA4 : rd_rsp_data <= 32'h000300A0;
                16'h0CBC : rd_rsp_data <= 32'h28000000;
                16'h0CD8 : rd_rsp_data <= 32'h64B22427;
                16'h0CDC : rd_rsp_data <= 32'h00766932;
                16'h0CE0 : rd_rsp_data <= 32'h00222222;
                16'h0CE4 : rd_rsp_data <= 32'h00040000;
                16'h0CE8 : rd_rsp_data <= 32'h77644302;
                16'h0CEC : rd_rsp_data <= 32'h2F97D40C;
                16'h0CF0 : rd_rsp_data <= 32'h00C70000;
                16'h0CF4 : rd_rsp_data <= 32'h00230000;
                16'h0CFC : rd_rsp_data <= 32'h80000000;
                16'h0D00 : rd_rsp_data <= 32'h00080740;
                16'h0D04 : rd_rsp_data <= 32'h00020403;
                16'h0D08 : rd_rsp_data <= 32'h0000907F;
                16'h0D0C : rd_rsp_data <= 32'h20010201;
                16'h0D10 : rd_rsp_data <= 32'hA0633333;
                16'h0D14 : rd_rsp_data <= 32'h3333BC43;
                16'h0D18 : rd_rsp_data <= 32'h7A8F5B6B;
                16'h0D1C : rd_rsp_data <= 32'h0000007F;
                16'h0D2C : rd_rsp_data <= 32'hCC979975;
                16'h0D34 : rd_rsp_data <= 32'h40608000;
                16'h0D3C : rd_rsp_data <= 32'h00127353;
                16'h0D50 : rd_rsp_data <= 32'h6437140A;
                16'h0D58 : rd_rsp_data <= 32'h00000282;
                16'h0D5C : rd_rsp_data <= 32'h30032064;
                16'h0D60 : rd_rsp_data <= 32'h4653DA68;
                16'h0D64 : rd_rsp_data <= 32'h04518A3C;
                16'h0D68 : rd_rsp_data <= 32'h00002101;
                16'h0D6C : rd_rsp_data <= 32'h2A201C16;
                16'h0D70 : rd_rsp_data <= 32'h1812362E;
                16'h0D74 : rd_rsp_data <= 32'h322C2220;
                16'h0D78 : rd_rsp_data <= 32'h000E3C24;
                16'h0D80 : rd_rsp_data <= 32'h01081008;
                16'h0D84 : rd_rsp_data <= 32'h00000800;
                16'h0D88 : rd_rsp_data <= 32'hF0B50000;
                16'h0DA0 : rd_rsp_data <= 32'h054D0B85;
                16'h0DA4 : rd_rsp_data <= 32'h0034059D;
                16'h0DA8 : rd_rsp_data <= 32'h0000002B;
                16'h0DAC : rd_rsp_data <= 32'h07900790;
                16'h0DB0 : rd_rsp_data <= 32'h0B040CC6;
                16'h0DB4 : rd_rsp_data <= 32'h0B040CC6;
                16'h0DB8 : rd_rsp_data <= 32'h010B00D5;
                16'h0DBC : rd_rsp_data <= 32'h0B470AB4;
                16'h0DC4 : rd_rsp_data <= 32'h03FA0000;
                16'h0DC8 : rd_rsp_data <= 32'h00000018;
                16'h0DCC : rd_rsp_data <= 32'h00000002;
                16'h0DD0 : rd_rsp_data <= 32'h00001108;
                16'h0DD4 : rd_rsp_data <= 32'h00000007;
                16'h0DD8 : rd_rsp_data <= 32'h80E10823;
                16'h0DDC : rd_rsp_data <= 32'h80003102;
                16'h0DE0 : rd_rsp_data <= 32'h0CC60CC6;
                16'h0DE8 : rd_rsp_data <= 32'h0002447C;
                16'h0DF4 : rd_rsp_data <= 32'h205E7000;
                16'h0DF8 : rd_rsp_data <= 32'h00000028;
                16'h0E00 : rd_rsp_data <= 32'h29292929;
                16'h0E04 : rd_rsp_data <= 32'h29292929;
                16'h0E08 : rd_rsp_data <= 32'h03902330;
                16'h0E0C : rd_rsp_data <= 32'h00000007;
                16'h0E10 : rd_rsp_data <= 32'h2B2B2B2B;
                16'h0E14 : rd_rsp_data <= 32'h292B2B2B;
                16'h0E18 : rd_rsp_data <= 32'h29292929;
                16'h0E1C : rd_rsp_data <= 32'h27292929;
                16'h0E28 : rd_rsp_data <= 32'h00000058;
                16'h0E30 : rd_rsp_data <= 32'h01008C00;
                16'h0E34 : rd_rsp_data <= 32'h01008C00;
                16'h0E38 : rd_rsp_data <= 32'h821608FF;
                16'h0E3C : rd_rsp_data <= 32'h281608FF;
                16'h0E40 : rd_rsp_data <= 32'h81037C02;
                16'h0E44 : rd_rsp_data <= 32'h01004800;
                16'h0E48 : rd_rsp_data <= 32'hF8000000;
                16'h0E4C : rd_rsp_data <= 32'h0046A891;
                16'h0E50 : rd_rsp_data <= 32'h38008C1C;
                16'h0E54 : rd_rsp_data <= 32'h18008C1C;
                16'h0E58 : rd_rsp_data <= 32'h821608FF;
                16'h0E5C : rd_rsp_data <= 32'h281608FF;
                16'h0E60 : rd_rsp_data <= 32'h00000048;
                16'h0E68 : rd_rsp_data <= 32'h0FC05656;
                16'h0E6C : rd_rsp_data <= 32'h03C09696;
                16'h0E70 : rd_rsp_data <= 32'h03C09696;
                16'h0E74 : rd_rsp_data <= 32'h0C005656;
                16'h0E78 : rd_rsp_data <= 32'h0C005656;
                16'h0E7C : rd_rsp_data <= 32'h0C005656;
                16'h0E80 : rd_rsp_data <= 32'h0C005656;
                16'h0E84 : rd_rsp_data <= 32'h03C09696;
                16'h0E88 : rd_rsp_data <= 32'h0C005656;
                16'h0E8C : rd_rsp_data <= 32'h03C09696;
                16'h0E90 : rd_rsp_data <= 32'h000001EC;
                16'h0E94 : rd_rsp_data <= 32'h01000000;
                16'h0E98 : rd_rsp_data <= 32'h0000007C;
                16'h0EA0 : rd_rsp_data <= 32'h0012C088;
                16'h0EA4 : rd_rsp_data <= 32'h01080000;
                16'h0EA8 : rd_rsp_data <= 32'h00001330;
                16'h0EAC : rd_rsp_data <= 32'h27FBA000;
                16'h0EB0 : rd_rsp_data <= 32'h000003C4;
                16'h0EB4 : rd_rsp_data <= 32'h01030000;
                16'h0EB8 : rd_rsp_data <= 32'h00000078;
                16'h0EBC : rd_rsp_data <= 32'h00020000;
                16'h0EC0 : rd_rsp_data <= 32'h00056F28;
                16'h0EC4 : rd_rsp_data <= 32'h01050000;
                16'h0EC8 : rd_rsp_data <= 32'h00000AC0;
                16'h0ED0 : rd_rsp_data <= 32'h03C09696;
                16'h0ED4 : rd_rsp_data <= 32'h03C09696;
                16'h0ED8 : rd_rsp_data <= 32'h03C09696;
                16'h0EDC : rd_rsp_data <= 32'h0000D6D6;
                16'h0EE0 : rd_rsp_data <= 32'h0000D6D6;
                16'h0EE4 : rd_rsp_data <= 32'hB0000C1C;
                16'h0EE8 : rd_rsp_data <= 32'h00000001;
                16'h0EEC : rd_rsp_data <= 32'h0FC01616;
                16'h0EF0 : rd_rsp_data <= 32'h83040000;
                16'h0EF4 : rd_rsp_data <= 32'h00000003;
                16'h0F00 : rd_rsp_data <= 32'h00000300;
                16'h0F14 : rd_rsp_data <= 32'h00000003;
                16'h0F80 : rd_rsp_data <= 32'h00000003;
                16'h0F84 : rd_rsp_data <= 32'h00000008;
                16'h0F88 : rd_rsp_data <= 32'h00000025;
                16'h0F94 : rd_rsp_data <= 32'h01570000;
                16'h0FA0 : rd_rsp_data <= 32'h03AB0000;
                16'h0FA4 : rd_rsp_data <= 32'h00010E9F;
                16'h0FA8 : rd_rsp_data <= 32'h0000CA0D;
                16'h0FAC : rd_rsp_data <= 32'h0002DC0E;
                16'h0FB0 : rd_rsp_data <= 32'h0940040A;
                16'h0FB4 : rd_rsp_data <= 32'h000098B6;
                16'h2000 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2004 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2008 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h200C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2010 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2014 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2018 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h201C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2020 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2024 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2028 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h202C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2030 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2034 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2038 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h203C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2040 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2044 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2048 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h204C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2050 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2054 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2058 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h205C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2060 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2064 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2068 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h206C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2070 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2074 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2078 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h207C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2080 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2084 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2088 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h208C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2090 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2094 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2098 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h209C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h20FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2100 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2104 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2108 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h210C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2110 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2114 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2118 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h211C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2120 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2124 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2128 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h212C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2130 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2134 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2138 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h213C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2140 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2144 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2148 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h214C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2150 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2154 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2158 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h215C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2160 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2164 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2168 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h216C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2170 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2174 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2178 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h217C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2180 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2184 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2188 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h218C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2190 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2194 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2198 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h219C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h21FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2200 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2204 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2208 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h220C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2210 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2214 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2218 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h221C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2220 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2224 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2228 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h222C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2230 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2234 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2238 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h223C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2240 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2244 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2248 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h224C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2250 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2254 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2258 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h225C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2260 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2264 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2268 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h226C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2270 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2274 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2278 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h227C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2280 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2284 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2288 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h228C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2290 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2294 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2298 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h229C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h22FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2300 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2304 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2308 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h230C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2310 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2314 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2318 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h231C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2320 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2324 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2328 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h232C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2330 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2334 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2338 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h233C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2340 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2344 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2348 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h234C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2350 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2354 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2358 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h235C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2360 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2364 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2368 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h236C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2370 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2374 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2378 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h237C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2380 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2384 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2388 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h238C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2390 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2394 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2398 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h239C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h23FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2400 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2404 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2408 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h240C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2410 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2414 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2418 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h241C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2420 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2424 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2428 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h242C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2430 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2434 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2438 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h243C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2440 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2444 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2448 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h244C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2450 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2454 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2458 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h245C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2460 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2464 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2468 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h246C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2470 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2474 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2478 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h247C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2480 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2484 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2488 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h248C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2490 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2494 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2498 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h249C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h24FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2500 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2504 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2508 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h250C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2510 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2514 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2518 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h251C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2520 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2524 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2528 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h252C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2530 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2534 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2538 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h253C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2540 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2544 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2548 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h254C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2550 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2554 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2558 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h255C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2560 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2564 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2568 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h256C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2570 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2574 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2578 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h257C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2580 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2584 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2588 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h258C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2590 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2594 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2598 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h259C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h25FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2600 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2604 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2608 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h260C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2610 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2614 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2618 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h261C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2620 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2624 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2628 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h262C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2630 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2634 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2638 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h263C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2640 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2644 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2648 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h264C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2650 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2654 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2658 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h265C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2660 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2664 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2668 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h266C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2670 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2674 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2678 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h267C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2680 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2684 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2688 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h268C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2690 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2694 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2698 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h269C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h26FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2700 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2704 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2708 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h270C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2710 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2714 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2718 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h271C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2720 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2724 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2728 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h272C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2730 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2734 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2738 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h273C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2740 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2744 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2748 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h274C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2750 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2754 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2758 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h275C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2760 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2764 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2768 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h276C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2770 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2774 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2778 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h277C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2780 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2784 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2788 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h278C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2790 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2794 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2798 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h279C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h27FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2800 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2804 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2808 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h280C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2810 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2814 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2818 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h281C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2820 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2824 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2828 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h282C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2830 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2834 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2838 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h283C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2840 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2844 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2848 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h284C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2850 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2854 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2858 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h285C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2860 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2864 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2868 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h286C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2870 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2874 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2878 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h287C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2880 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2884 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2888 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h288C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2890 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2894 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2898 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h289C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h28FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2900 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2904 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2908 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h290C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2910 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2914 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2918 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h291C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2920 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2924 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2928 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h292C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2930 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2934 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2938 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h293C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2940 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2944 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2948 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h294C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2950 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2954 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2958 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h295C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2960 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2964 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2968 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h296C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2970 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2974 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2978 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h297C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2980 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2984 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2988 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h298C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2990 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2994 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2998 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h299C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h29FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2A9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ABC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ACC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ADC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2AFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2B9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2BFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2C9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2CFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2D9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2DFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2E9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ECC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ED0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ED4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2ED8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2EFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2F9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h2FFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3000 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3004 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3008 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h300C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3010 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3014 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3018 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h301C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3020 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3024 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3028 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h302C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3030 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3034 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3038 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h303C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3040 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3044 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3048 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h304C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3050 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3054 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3058 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h305C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3060 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3064 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3068 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h306C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3070 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3074 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3078 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h307C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3080 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3084 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3088 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h308C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3090 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3094 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3098 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h309C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h30FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3100 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3104 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3108 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h310C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3110 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3114 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3118 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h311C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3120 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3124 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3128 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h312C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3130 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3134 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3138 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h313C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3140 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3144 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3148 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h314C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3150 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3154 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3158 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h315C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3160 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3164 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3168 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h316C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3170 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3174 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3178 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h317C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3180 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3184 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3188 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h318C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3190 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3194 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3198 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h319C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h31FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3200 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3204 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3208 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h320C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3210 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3214 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3218 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h321C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3220 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3224 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3228 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h322C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3230 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3234 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3238 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h323C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3240 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3244 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3248 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h324C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3250 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3254 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3258 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h325C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3260 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3264 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3268 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h326C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3270 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3274 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3278 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h327C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3280 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3284 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3288 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h328C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3290 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3294 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3298 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h329C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h32FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3300 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3304 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3308 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h330C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3310 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3314 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3318 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h331C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3320 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3324 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3328 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h332C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3330 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3334 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3338 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h333C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3340 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3344 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3348 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h334C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3350 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3354 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3358 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h335C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3360 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3364 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3368 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h336C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3370 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3374 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3378 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h337C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3380 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3384 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3388 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h338C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3390 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3394 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3398 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h339C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h33FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3400 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3404 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3408 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h340C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3410 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3414 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3418 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h341C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3420 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3424 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3428 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h342C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3430 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3434 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3438 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h343C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3440 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3444 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3448 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h344C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3450 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3454 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3458 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h345C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3460 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3464 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3468 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h346C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3470 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3474 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3478 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h347C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3480 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3484 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3488 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h348C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3490 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3494 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3498 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h349C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h34FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3500 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3504 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3508 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h350C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3510 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3514 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3518 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h351C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3520 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3524 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3528 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h352C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3530 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3534 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3538 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h353C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3540 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3544 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3548 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h354C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3550 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3554 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3558 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h355C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3560 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3564 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3568 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h356C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3570 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3574 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3578 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h357C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3580 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3584 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3588 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h358C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3590 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3594 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3598 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h359C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h35FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3600 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3604 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3608 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h360C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3610 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3614 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3618 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h361C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3620 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3624 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3628 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h362C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3630 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3634 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3638 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h363C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3640 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3644 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3648 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h364C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3650 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3654 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3658 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h365C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3660 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3664 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3668 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h366C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3670 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3674 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3678 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h367C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3680 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3684 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3688 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h368C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3690 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3694 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3698 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h369C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h36FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3700 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3704 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3708 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h370C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3710 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3714 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3718 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h371C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3720 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3724 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3728 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h372C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3730 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3734 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3738 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h373C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3740 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3744 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3748 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h374C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3750 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3754 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3758 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h375C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3760 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3764 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3768 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h376C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3770 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3774 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3778 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h377C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3780 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3784 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3788 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h378C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3790 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3794 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3798 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h379C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h37FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3800 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3804 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3808 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h380C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3810 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3814 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3818 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h381C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3820 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3824 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3828 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h382C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3830 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3834 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3838 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h383C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3840 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3844 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3848 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h384C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3850 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3854 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3858 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h385C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3860 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3864 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3868 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h386C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3870 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3874 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3878 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h387C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3880 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3884 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3888 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h388C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3890 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3894 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3898 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h389C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h38FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3900 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3904 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3908 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h390C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3910 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3914 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3918 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h391C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3920 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3924 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3928 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h392C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3930 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3934 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3938 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h393C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3940 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3944 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3948 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h394C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3950 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3954 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3958 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h395C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3960 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3964 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3968 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h396C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3970 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3974 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3978 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h397C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3980 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3984 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3988 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h398C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3990 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3994 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3998 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h399C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39A0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39A4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39A8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39AC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39B0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39B4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39B8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39BC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39C0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39C4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39C8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39CC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39D0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39D4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39D8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39DC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39E0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39E4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39E8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39EC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39F0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39F4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39F8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h39FC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3A9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ABC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ACC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ADC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3AFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3B9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3BFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3C9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3CFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3D9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3DFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3E9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ECC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ED0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ED4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3ED8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3EFC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F00 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F04 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F08 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F0C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F10 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F14 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F18 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F1C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F20 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F24 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F28 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F2C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F30 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F34 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F38 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F3C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F40 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F44 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F48 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F4C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F50 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F54 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F58 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F5C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F60 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F64 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F68 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F6C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F70 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F74 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F78 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F7C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F80 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F84 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F88 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F8C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F90 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F94 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F98 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3F9C : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FA0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FA4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FA8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FAC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FB0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FB4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FB8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FBC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FC0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FC4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FC8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FCC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FD0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FD4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FD8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FDC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FE0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FE4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FE8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FEC : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FF0 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FF4 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FF8 : rd_rsp_data <= 32'hEAEAEAEA;
                16'h3FFC : rd_rsp_data <= 32'hEAEAEAEA;
                default: rd_rsp_data <= 32'h00000000;
            endcase
        end else if (dwr_valid) begin
            case (({dwr_addr[31:24], dwr_addr[23:16], dwr_addr[15:08], dwr_addr[07:00]} - (base_address_register & 32'hFFFFFFF0)) & 32'hFFFF)
                //Dont be scared
            endcase
        end else begin
            rd_rsp_data <= 32'h00000000;
        end
    end
            
endmodule
